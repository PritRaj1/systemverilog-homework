`include "util.svh"

module testbench;

  logic [3:0] d0, d1, d2, d3;
  logic [1:0] sel;
  logic [3:0] y;

  mux_4_1 inst (
      .d0 (d0),
      .d1 (d1),
      .d2 (d2),
      .d3 (d3),
      .sel(sel),
      .y  (y)
  );

  task test(input [3:0] td0, td1, td2, td3, input [1:0] tsel, input [3:0] ty);

    {d0, d1, d2, d3, sel} = {td0, td1, td2, td3, tsel};

    #1;

    if (y !== ty) begin
      $display("FAIL %s", `__FILE__);
      $display("++ INPUT    => {%s, %s, %s, %s, %s}", `PH(d0), `PH(d1), `PH(d2), `PH(d3), `PH(sel));
      $display("++ EXPECTED => {%s}", `PH(ty));
      $display("++ ACTUAL   => {%s}", `PH(y));
      $finish(1);
    end

  endtask

  initial begin
    test('ha, 'hb, 'hc, 'hd, 0, 'ha);
    test('ha, 'hb, 'hc, 'hd, 1, 'hb);
    test('ha, 'hb, 'hc, 'hd, 2, 'hc);
    test('ha, 'hb, 'hc, 'hd, 3, 'hd);

    test(7, 10, 3, 'x, 0, 7);
    test(7, 10, 3, 'x, 1, 10);
    test(7, 10, 3, 'x, 2, 3);
    test(7, 10, 3, 'x, 3, 'x);

    $display("PASS %s", `__FILE__);
    $finish;
  end

endmodule
